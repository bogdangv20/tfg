-- DDR controller
  constant CFG_DDR2SP  		   : integer := CONFIG_DDR2SP;
  constant CFG_DDR2SP_INIT  	   : integer := CONFIG_DDR2SP_INIT;
  constant CFG_DDR2SP_FREQ   	   : integer := CONFIG_DDR2SP_FREQ;
  constant CFG_DDR2SP_TRFC   	   : integer := CONFIG_DDR2SP_TRFC;
  constant CFG_DDR2SP_DATAWIDTH    : integer := CONFIG_DDR2SP_DATAWIDTH;
  constant CFG_DDR2SP_FTEN         : integer := CONFIG_DDR2SP_FTEN;
  constant CFG_DDR2SP_FTWIDTH      : integer := CONFIG_DDR2SP_FTWIDTH;
  constant CFG_DDR2SP_COL    	   : integer := CONFIG_DDR2SP_COL;
  constant CFG_DDR2SP_SIZE  	   : integer := CONFIG_DDR2SP_MBYTE;
  constant CFG_DDR2SP_DELAY0 	   : integer := CONFIG_DDR2SP_DELAY0;
  constant CFG_DDR2SP_DELAY1 	   : integer := CONFIG_DDR2SP_DELAY1;
  constant CFG_DDR2SP_DELAY2 	   : integer := CONFIG_DDR2SP_DELAY2;
  constant CFG_DDR2SP_DELAY3 	   : integer := CONFIG_DDR2SP_DELAY3;
  constant CFG_DDR2SP_DELAY4 	   : integer := CONFIG_DDR2SP_DELAY4;
  constant CFG_DDR2SP_DELAY5 	   : integer := CONFIG_DDR2SP_DELAY5;
  constant CFG_DDR2SP_DELAY6 	   : integer := CONFIG_DDR2SP_DELAY6;
  constant CFG_DDR2SP_DELAY7 	   : integer := CONFIG_DDR2SP_DELAY7;
  constant CFG_DDR2SP_NOSYNC       : integer := CONFIG_DDR2SP_NOSYNC;
  constant CFG_DDR2SP_OBFUSCATION : integer := CONFIG_DDR2SP_OBFUSCATION;
  constant CFG_DDR2SP_OBFUSCATION_START : integer := 16#CONFIG_DDR2SP_OBFUSCATION_START#;
  constant CFG_DDR2SP_OBFUSCATION_END : integer := 16#CONFIG_DDR2SP_OBFUSCATION_END#;
